module addr_gen
(
 input wire[31:0] address_in,
 output wire [31:0] address_out
 );
 
	 assign address_out = address_in ;


endmodule