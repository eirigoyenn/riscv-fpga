module sum4
(
 input wire[31:0] val_in,
 output wire [31:0] val_out
 );
 
	 assign val_out = val_in + 4;


endmodule